////////////////////////////////////////////////////////////////////////////////
// SubModule BLE
// Created   2/25/2017 3:22:46 PM
////////////////////////////////////////////////////////////////////////////////

module BLE (O\C\P\, Antenna, RXD, TXD);

input  O\C\P\;
inout  Antenna;
inout  RXD;
inout  TXD;


endmodule
////////////////////////////////////////////////////////////////////////////////
